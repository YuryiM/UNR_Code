library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package fsm_types is
    type state_type is (Reset, A, B, C, D, E, F, G, H, I, J, K);
end fsm_types;